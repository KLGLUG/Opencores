module main;
	initial
		begin
			$display("This is the first verilog code");
			$finish ;
		end
endmodule
